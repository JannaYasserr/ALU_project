module comp_tb;
reg [7:0] A, B;
wire E,G,L;

comp_beh uut(A, B, E,G,L);

initial 
begin

A=8'b00011100;
B=8'b00010100;

#100;
A=8'b01111100;
B=8'b00010100;

#100;
A=8'b10011100;
B=8'b00010100;

#100;
A=8'b10011100;
B=8'b10010100;

#100;
A=8'b00011100;
B=8'b00011100;

#100;
A=8'b11011100;
B=8'b11010100;

#100;
A=8'b00000100;
B=8'b00010100;

#100;

end
endmodule
