module and_struct(A,B,S);
input [7:0] A,B;
output [7:0] S;


and a1(S[0],A[0],B[0]);
and a2(S[1],A[1],B[1]);
and a3(S[2],A[2],B[2]);
and a4(S[3],A[3],B[3]);
and a5(S[4],A[4],B[4]);
and a6(S[5],A[5],B[5]);
and a7(S[6],A[6],B[6]);
and a8(S[7],A[7],B[7]);

endmodule
