module comp_beh(A,B,E,G,L);
input [7:0] A , B;
output reg E,G,L;
always @(*)
if ((A[7]<B[7])|((A[7]==B[7])&(A[6]>B[6]))|((A[7]==B[7])&(A[6]==B[6])&(A[5]>B[5]))|((A[7]==B[7])&(A[6]==B[6])&(A[5]==B[5])&(A[4]>B[4]))|((A[7]==B[7])&(A[6]==B[6])&(A[5]==B[5])&(A[4]==B[4])&(A[3]>B[3]))|((A[7]==B[7])&(A[6]==B[6])&(A[5]==B[5])&(A[4]==B[4])&(A[3]==B[3])&(A[2]>B[2]))|((A[7]==B[7])&(A[6]==B[6])&(A[5]==B[5])&(A[4]==B[4])&(A[3]==B[3])&(A[2]==B[2])&(A[1]>B[1]))|((A[7]==B[7])&(A[6]==B[6])&(A[5]==B[5])&(A[4]==B[4])&(A[3]==B[3])&(A[2]==B[2])&(A[1]==B[1])&(A[0]>B[0])))
begin
G=1;
L=0;
E=0;
end
else if((A[7]==B[7])&(A[6]==B[6])&(A[5]==B[5])&(A[4]==B[4])&(A[3]==B[3])&(A[2]==B[2])&(A[1]==B[1])&(A[0]==B[0]))
begin
G=0;
L=0;
E=1;
end
else
begin
G=0;
L=1;
E=0;
end

endmodule
