module topAU_tb;
reg [7:0] A,B;
reg S3,S2;
wire C,O,Z,E,G,L;
wire [7:0] S;

topAU uut(A,B,S3,S2,S,C,O,Z,E,G,L);

initial 
begin

A=8'b00011100;
B=8'b00010100;
S3=0;
S2=0;

#100;
A=8'b01111100;
B=8'b00010100;
S3=1;
S2=1;
#100;
A=8'b10011100;
B=8'b00010100;
S3=1;
S2=0;
#100;
A=8'b10011100;
B=8'b10010100;
S3=0;
S2=0;
#100;
A=8'b00011100;
B=8'b00011100;
S3=1;
S2=0;
#100;
A=8'b11011100;
B=8'b11010100;
S3=1;
S2=0;
#100;
A=8'b00000100;
B=8'b00010100;
S3=1;
S2=1;
#100;

end
endmodule
